LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ProgramCounter IS
	PORT (
		CLOCK : IN STD_LOGIC;
		PC_INC : IN STD_LOGIC_VECTOR(0 TO 31);
		PC : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"
	);
END ProgramCounter;

ARCHITECTURE PC OF ProgramCounter IS
BEGIN
	PROCESS (CLOCK, PC_INC)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN
			PC <= PC_INC;
		END IF;
	END PROCESS;
END;