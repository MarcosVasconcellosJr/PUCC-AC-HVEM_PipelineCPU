LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

-- This component implements a pipeline register, in this case (is the) first register of the first stage
ENTITY Reg_Pipe_IFID IS
	PORT (
		-- IN --
		CLOCK : IN STD_LOGIC;
		IN_PC_MAIS_4 : IN STD_LOGIC_VECTOR(0 TO 31); -- PC Increment
		IN_INSTR_MEM : IN STD_LOGIC_VECTOR(0 TO 31); -- Instruction
		-- OUT --
		OUT_PC_MAIS_4 : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"; -- Out PC Increment
		OUT_INSTR_MEM : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"); -- Out instruction
END Reg_Pipe_IFID;

ARCHITECTURE REG_PIPE OF Reg_Pipe_IFID IS
BEGIN
	PROCESS (CLOCK)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN
			OUT_INSTR_MEM <= IN_INSTR_MEM;
			OUT_PC_MAIS_4 <= IN_PC_MAIS_4;
		END IF;
	END PROCESS;
END;