LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Cpu IS
    GENERIC (DATA_SIZE : INTEGER := 32); -- Generic data size to map in components
    PORT (
        CLOCK : IN STD_LOGIC
    );
END Cpu;

ARCHITECTURE CPU OF Cpu IS

    -- Control Unit - PORT MAP
    COMPONENT ControlUnit
        PORT (
            WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            EX : OUT STD_LOGIC_VECTOR(0 TO 4);
            SIGNAL_JUMP : OUT STD_LOGIC_VECTOR(0 TO 1);
            OP_CODE : IN STD_LOGIC_VECTOR(0 TO 5)
        );
    END COMPONENT;

    -- ShiftLeft - PORT MAP
    COMPONENT ShiftLeft
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 31);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- ShiftLeft2_26to28 - PORT MAP
    COMPONENT ShiftLeft2_26to28
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 25);
            X : OUT STD_LOGIC_VECTOR(0 TO 27)
        );
    END COMPONENT;

    -- Signal Extend - PORT MAP
    COMPONENT SignalExtend
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 15);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- Generic2to1Mux - PORT MAP
    COMPONENT Generic2to1Mux
        PORT (
            CONTROL : IN STD_LOGIC;
            A : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
            B : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);

            X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1)
        );
    END COMPONENT;

    --  Generic3to1Mux - PORT MAP
    COMPONENT Generic3to1Mux
        PORT (
            JUMP_SIGNAL : IN STD_LOGIC_VECTOR (0 TO 1);
            A, B, C : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);

            X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1)
        );
    END COMPONENT;

    -- Alu - PORT MAP
    COMPONENT Alu
        PORT (
            RS_DATA : IN STD_LOGIC_VECTOR(0 TO 31);
            RT_DATA : IN STD_LOGIC_VECTOR(0 TO 31);
            ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1);

            ALU_OUT : OUT STD_LOGIC_VECTOR(0 TO 31);
            ZERO : OUT STD_LOGIC
        );
    END COMPONENT;

    -- Data Memory - PORT MAP
    COMPONENT DataMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
            CLOCK : IN STD_LOGIC;
            MEM_WRITE : IN STD_LOGIC;
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 31);
            MEM_READ : IN STD_LOGIC;

            READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- InstructionMemory - PORT MAP
    COMPONENT InstructionMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
            INSTRUCTION : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"
        );
    END COMPONENT;

    -- PCIncrement - PORT MAP
    COMPONENT PCIncrement
        PORT (
            PC : IN STD_LOGIC_VECTOR (0 TO 31);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- Reg_Pipe_IFID - PORT MAP
    COMPONENT Reg_Pipe_IFID
        PORT (
            IN_PC_MAIS_4 : IN STD_LOGIC_VECTOR(0 TO 31);
            IN_INSTR_MEM : IN STD_LOGIC_VECTOR(0 TO 31);
            IN_PC_WRITE : IN STD_LOGIC_VECTOR;

            OUT_PC_MAIS_4 : OUT STD_LOGIC_VECTOR(0 TO 31);
            OUT_INSTR_MEM : OUT STD_LOGIC_VECTOR(0 TO 31);
            OUT_PC_WRITE : OUT STD_LOGIC_VECTOR
        );
    END COMPONENT;

    -- Reg_Pipe_IDEX - PORT MAP
    COMPONENT Reg_Pipe_IDEX
        PORT (
            CLOCK : IN STD_LOGIC;
            IDEX_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            IDEX_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            IDEX_IN_EX : IN STD_LOGIC_VECTOR(0 TO 4);
            IDEX_IN_PC : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_READ1 : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_IMED : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_RT : IN STD_LOGIC_VECTOR(0 TO 4);
            IDEX_IN_RD : IN STD_LOGIC_VECTOR(0 TO 4);
            IN_PC_WRITE : IN STD_LOGIC_VECTOR;

            IDEX_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            IDEX_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            IDEX_OUT_EX : OUT STD_LOGIC_VECTOR(0 TO 4);
            IDEX_OUT_PC : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_READ1 : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_IMED : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_RT : OUT STD_LOGIC_VECTOR(0 TO 4);
            IDEX_OUT_RD : OUT STD_LOGIC_VECTOR(0 TO 4);
            OUT_PC_WRITE : OUT STD_LOGIC_VECTOR
        );
    END COMPONENT;

    -- Reg_Pipe_EXMEM - PORT MAP
    COMPONENT Reg_Pipe_EXMEM
        PORT (
            CLOCK : IN STD_LOGIC;
            EXMEM_IN_ZERO : IN STD_LOGIC;
            EXMEM_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_IN_RESULT_ADDER : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 4);
            IN_PC_WRITE : IN STD_LOGIC_VECTOR;

            EXMEM_OUT_ZERO : OUT STD_LOGIC;
            EXMEM_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_OUT_RESULT_ADDER : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 4);
            OUT_PC_WRITE : OUT STD_LOGIC_VECTOR
        );
    END COMPONENT;

    -- Reg_Pipe_MEMWB - PORT MAP
    COMPONENT Reg_Pipe_MEMWB
        PORT (
            CLOCK : IN STD_LOGIC;
            MEMWB_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 31);
            MEMWB_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 4);
            MEMWB_IN_READ_DATA : IN STD_LOGIC_VECTOR(0 TO 31);

            MEMWB_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
            MEMWB_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 4);
            MEMWB_OUT_READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- FileRegister - PORT MAP
    COMPONENT FileRegister
        PORT (
            REGWRITE : IN STD_LOGIC;
            CLOCK : IN STD_LOGIC;
            READ_REGISTER_1 : IN STD_LOGIC_VECTOR(0 TO 4);
            READ_REGISTER_2 : IN STD_LOGIC_VECTOR(0 TO 4);
            WRITE_REGISTER : IN STD_LOGIC_VECTOR(0 TO 4);
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 31);

            READ_DATA_1 : OUT STD_LOGIC_VECTOR(0 TO 31);
            READ_DATA_2 : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    --******************** INSTRUCTION FETCH ********************--

    -- SIGNALS - TO CONTROL COMPONENT INTERACTION IN EXECUTION TIME
    SIGNAL SIG_PC_SRC : STD_LOGIC;
    SIGNAL SIG_JUMP : STD_LOGIC;

    -- WIRES - TO CONNECT PORT MAP BETWEEN COMPONENTS
    SIGNAL WIRE_OUT_PC_INC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_PC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_PC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_JUMP : STD_LOGIC_VECTOR(0 TO 31); --Used to connect mux 
    SIGNAL WIRE_INST_MEM_IFID : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_PC : STD_LOGIC_VECTOR(0 TO 31);

    --******************** COMPONENTS INSTRUCTION FETCH ********************--

    INST_MEM : InstructionMemory PORT MAP(WIRE_PC_INST_MEM, WIRE_INST_MEM_IFID);
    PC_INC : PCIncrement PORT MAP(WIRE_OUT_PC, WIRE_OUT_PC_INC);
    PC : ProgramCounter PORT MAP(CLOCK, WIRE_OUT_PC_INC, WIRE_PC);
    MUX_PC : Generic2to1Mux PORT MAP(TODO : AQUI O QUE VIER DO BRANCH, WIRE_OUT_PC_INC);

    --******************** REG_PIPELINE IF/ID ********************--

    IFID : Pipe_Reg_IFID
    PORT MAP(
        -- IN
        WIRE_OUT_PC_INC, WIRE_INST_MEM_IFID,
        -- OUT
        WIRE_PC_INC_IFID_TO_IDEX, WIRE_OUT_IFID_INSTRUCTION
    );

    --******************** SIGNALS AND WIRES OF INSTRUCTION DECODE STAGE     ********************--

    --WIRES
    SIGNAL WIRE_PC_INC_IFID_TO_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_IFID_INSTRUCTION : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_READ_DATA1_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_READ_DATA2_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_SIGNAL_EXTEND_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    -- Control Unit
    SIGNAL WIRE_UC_IDEX_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_UC_IDEX_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_UC_IDEX_EX : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_UC_JUMP_SIGNAL : STD_LOGIC_VECTOR(0 TO 1); --TODO TROCAR NOME

    SIGNAL WIRE_IDEX_WB_EXMEM_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_IDEX_MEM_EXMEM_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_PC_INC_IDEX_TO_ADDER : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_READ1_ALU_A : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_READ2_MUX_ALU_B : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_IDEX_IMED : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_RT_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_RD_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 31);

    --******************** COMPONENTS INSTRUCTION DECODE     ********************--

    FILE_REG : FileRegister PORT MAP(TODO : REGWRITE, CLOCK, WIRE_OUT_IFID_INSTRUCTION(6 TO 11), WIRE_OUT_IFID_INSTRUCTION(12 TO 16), TODO : WRITE_REGISTER, TODO : WRITEDATA VEM DO MUX WB, WIRE_READ_DATA1_IDEX, WIRE_READ_DATA2_IDEX);
    SIGNAL_EXTEND : SignExtend PORT MAP(WIRE_OUT_IFID_INSTRUCTION(0 TO 15), WIRE_SIGNAL_EXTEND_IDEX);
    UC : ControlUnit PORT MAP(WIRE_UC_IDEX_WB, WIRE_UC_IDEX_MEM, WIRE_UC_IDEX_EX, WIRE_UC_JUMP_SIGNAL, WIRE_OUT_IFID_INSTRUCTION(0 TO 5));

    --******************** REG_PIPELINE ID/EX ********************--

    IDEX : Pipe_Reg_IDEX
    PORT MAP(
        -- IN
        CLOCK,
        WIRE_UC_IDEX_WB,
        WIRE_UC_IDEX_MEM,
        WIRE_UC_IDEX_EX,
        WIRE_PC_INC_IFID_TO_IDEX,
        WIRE_READ_DATA1_IDEX,
        WIRE_READ_DATA2_IDEX,
        WIRE_SIGNAL_EXTEND_IDEX,
        WIRE_OUT_IFID_INSTRUCTION(11 TO 15),
        WIRE_OUT_IFID_INSTRUCTION(16 TO 20),
        -- OUT
        WIRE_IDEX_WB_EXMEM_WB,
        WIRE_IDEX_MEM_EXMEM_MEM,
        WIRE_OUT_IDEX_EX,
        WIRE_PC_INC_IDEX_TO_ADDER,
        WIRE_IDEX_READ1_ALU_A,
        WIRE_IDEX_READ2_MUX_ALU_B,
        WIRE_OUT_IDEX_IMED,
        WIRE_IDEX_RT_MUX_REGDST,
        WIRE_IDEX_RD_MUX_REGDST
    );

    EXMEM : Pipe_Reg_EXMEM
    PORT MAP(
        -- IN
        CLOCK,
        WIRE_ALU_ZERO
        -- OUT
    );

    --******************** INSTRUCTION EXECUTION STAGE  ********************--
    
    --******************** COMPONENTS I NSTRUCTION EXECUTION  ********************--
    --******************** REG_PIPELINE EX/MEM ********************--

    --******************** SIGNALS AND WIRES OF INSTRUCTION MEMORY STAGE     ********************--
    --******************** COMPONENTS INSTRUCTION MEMORY     ********************--
    --******************** REG_PIPELINE EX/MEM ********************--

    --******************** SIGNALS AND WIRES OF INSTRUCTION WRITE BACK STAGE ********************--
    --******************** COMPONENTS INSTRUCTION WRITE BACK ********************--
    --******************** REG_PIPELINE EX/MEM ********************--

END;