LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FileRegister IS
    PORT (
        REGWRITE : IN STD_LOGIC;
        CLOCK : IN STD_LOGIC;
        READ_REGISTER_1 : IN STD_LOGIC_VECTOR(0 TO 4);
        READ_REGISTER_2 : IN STD_LOGIC_VECTOR(0 TO 4);
        WRITE_REGISTER : IN STD_LOGIC_VECTOR(0 TO 4);
        WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 31);
        READ_DATA_1 : OUT STD_LOGIC_VECTOR(0 TO 31);
        READ_DATA_2 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_REGS : OUT STD_LOGIC_VECTOR(0 TO 31)
    );
END FileRegister;

ARCHITECTURE REGS OF FileRegister IS
    TYPE REGISTER_TYPE IS ARRAY(0 TO 31) OF STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL REGISTERS : REGISTER_TYPE;
BEGIN
    PROCESS (CLOCK)
    BEGIN
        IF (CLOCK'EVENT AND CLOCK = '1' AND REGWRITE = '1' AND NOT (WRITE_REGISTER = "00000")) THEN
            REGISTERS(TO_INTEGER(UNSIGNED(WRITE_REGISTER))) <= WRITE_DATA;
        END IF;
    END PROCESS;

    DEB_REGS <= REGISTERS(TO_INTEGER(UNSIGNED(00010)));
    READ_DATA_1 <= REGISTERS(TO_INTEGER(UNSIGNED(READ_REGISTER_1)));
    READ_DATA_2 <= REGISTERS(TO_INTEGER(UNSIGNED(READ_REGISTER_2)));
END;