LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Reg_Pipe_EXMEM IS
    PORT (
        -- IN --
        CLOCK : IN STD_LOGIC;
        EXMEM_IN_ZERO : IN STD_LOGIC; -- ALU RESULTS EQUALS TO ZERO SIGNAL
        EXMEM_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1); -- POSITION: (0 - RegWrite, 1 - MEMtoREG)
        EXMEM_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2); -- POSITION: (0 - BRANCH, 1- MEMRead, 2 - MEMWrite)
        EXMEM_IN_RESULT_ADDER : IN STD_LOGIC_VECTOR(0 TO 31); -- ADDER RESULT
        EXMEM_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 31); -- ALU RESULT
        EXMEM_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 31); -- READ
        EXMEM_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 4); -- EXIT MUX, RT OR RD
        -- OUT --
        EXMEM_OUT_ZERO : OUT STD_LOGIC;
        EXMEM_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
        EXMEM_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
        EXMEM_OUT_RESULT_ADDER : OUT STD_LOGIC_VECTOR(0 TO 31);
        EXMEM_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
        EXMEM_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 31);
        EXMEM_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 4));
END Reg_Pipe_EXMEM;

ARCHITECTURE REG_PIPE OF Reg_Pipe_EXMEM IS

BEGIN
    PROCESS (CLOCK)
    BEGIN
        IF (CLOCK'EVENT AND CLOCK = '1') THEN
            EXMEM_OUT_ZERO <= EXMEM_IN_ZERO;
            EXMEM_OUT_WB <= EXMEM_IN_WB;
            EXMEM_OUT_MEM <= EXMEM_IN_MEM;
            EXMEM_OUT_RESULT_ADDER <= EXMEM_IN_RESULT_ADDER;
            EXMEM_OUT_RESULT_ULA <= EXMEM_IN_RESULT_ULA;
            EXMEM_OUT_READ2 <= EXMEM_IN_READ2;
            EXMEM_OUT_REGDST <= EXMEM_IN_REGDST;
        END IF;
    END PROCESS;
END REG_PIPE;