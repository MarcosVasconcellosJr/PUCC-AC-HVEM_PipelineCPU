LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ALU IS
	PORT (
		RS_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- REGISTER
		RT_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- REGISTER
		ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1); -- CODE OF THE ARITHMETIC OPERATION OPTION
		ALU_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0); -- WHERE WE WILL STORE THE RESULT OF THE ARITHMETIC OPERATION
		ZERO: OUT STD_LOGIC);
END ALU;

ARCHITECTURE ALU OF ALU IS
	SIGNAL AUX: STD_LOGIC_VECTOR(0 to 31);
BEGIN
	PROCESS (RS_DATA, RS_DATA, ALU_CODE)
	BEGIN
		-- SWITCH CASE TO DO THE RIGHT OPERATION BASED IN ALU_CODE
		CASE ALU_CODE IS
			WHEN "00" => AUX <= RS_DATA + RT_DATA;
			WHEN "01" => AUX <= RS_DATA - RT_DATA;
			WHEN "10" => AUX <= RS_DATA AND RT_DATA;
			WHEN "11" => AUX <= RS_DATA OR RT_DATA;
			WHEN OTHERS => AUX <= "00000000000000000000000000000000";
		END CASE;
				IF(AUX = "00000000000000000000000000000000") THEN
			ZERO <= '1';
		ELSE
			ZERO <= '0';
		END IF;
		
		ALU_OUT <= AUX;
	END PROCESS;
END ALU;