LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY InstructionMemory IS

    PORT (
        ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
        INSTRUCTION : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"
        );

END InstructionMemory;

ARCHITECTURE MEM OF InstructionMemory IS
    TYPE MEM_TYPE IS ARRAY(0 TO 400) OF STD_LOGIC_VECTOR(0 TO 7);
    SIGNAL MEMORY : MEM_TYPE;
BEGIN

    MEMORY(000) <= "00001000";
    MEMORY(001) <= "00100010";
    MEMORY(002) <= "00000000";
    MEMORY(003) <= "00001000";--addi $2,$1, 8 |=>  $2 = 8

    MEMORY(004) <= "00001100";
    MEMORY(005) <= "01000001";
    MEMORY(006) <= "00000000";
    MEMORY(007) <= "00000001";--subi $1, $2, 1 |=>  $1 = 8, $2 = 7

    MEMORY(008) <= "00000000";
    MEMORY(009) <= "00000000";
    MEMORY(010) <= "00000000";
    MEMORY(011) <= "00000000";

    MEMORY(012) <= "00000000";
    MEMORY(013) <= "00000000";
    MEMORY(014) <= "00000000";
    MEMORY(015) <= "00000000";

    MEMORY(016) <= "00000000";
    MEMORY(017) <= "00000000";
    MEMORY(018) <= "00000000";
    MEMORY(019) <= "00000000";

    MEMORY(020) <= "00000000";
    MEMORY(021) <= "00000000";
    MEMORY(022) <= "00000000";
    MEMORY(023) <= "00000000";

    MEMORY(024) <= "00000000";
    MEMORY(025) <= "00000000";
    MEMORY(026) <= "00000000";
    MEMORY(027) <= "00000000";

    MEMORY(028) <= "00000000";
    MEMORY(029) <= "00000000";
    MEMORY(030) <= "00000000";
    MEMORY(031) <= "00000000";

    MEMORY(032) <= "00000000";
    MEMORY(033) <= "00000000";
    MEMORY(034) <= "00000000";
    MEMORY(035) <= "00000000";

    MEMORY(036) <= "00000000";
    MEMORY(037) <= "00000000";
    MEMORY(038) <= "00000000";
    MEMORY(039) <= "00000000";

    MEMORY(040) <= "00000000";
    MEMORY(041) <= "00000000";
    MEMORY(042) <= "00000000";
    MEMORY(043) <= "00000000";

    MEMORY(044) <= "00000000";
    MEMORY(045) <= "00000000";
    MEMORY(046) <= "00000000";
    MEMORY(047) <= "00000000";

    MEMORY(048) <= "00000000";
    MEMORY(049) <= "00000000";
    MEMORY(050) <= "00000000";
    MEMORY(051) <= "00000000";

    MEMORY(052) <= "00000000";
    MEMORY(053) <= "00000000";
    MEMORY(054) <= "00000000";
    MEMORY(055) <= "00000000";

    MEMORY(056) <= "00000000";
    MEMORY(057) <= "00000000";
    MEMORY(058) <= "00000000";
    MEMORY(059) <= "00000000";

    MEMORY(060) <= "00000000";
    MEMORY(061) <= "00000000";
    MEMORY(062) <= "00000000";
    MEMORY(063) <= "00000000";

    MEMORY(064) <= "00000000";
    MEMORY(065) <= "00000000";
    MEMORY(066) <= "00000000";
    MEMORY(067) <= "00000000";

    MEMORY(068) <= "00000000";
    MEMORY(069) <= "00000000";
    MEMORY(070) <= "00000000";
    MEMORY(071) <= "00000000";

    MEMORY(072) <= "00000000";
    MEMORY(073) <= "00000000";
    MEMORY(074) <= "00000000";
    MEMORY(075) <= "00000000";

    MEMORY(076) <= "00000000";
    MEMORY(077) <= "00000000";
    MEMORY(078) <= "00000000";
    MEMORY(079) <= "00000000";

    MEMORY(080) <= "00000000";
    MEMORY(081) <= "00000000";
    MEMORY(082) <= "00000000";
    MEMORY(083) <= "00000000";

    MEMORY(084) <= "00000000";
    MEMORY(085) <= "00000000";
    MEMORY(086) <= "00000000";
    MEMORY(087) <= "00000000";

    MEMORY(088) <= "00000000";
    MEMORY(089) <= "00000000";
    MEMORY(090) <= "00000000";
    MEMORY(091) <= "00000000";

    MEMORY(092) <= "00000000";
    MEMORY(093) <= "00000000";
    MEMORY(094) <= "00000000";
    MEMORY(095) <= "00000000";

    MEMORY(096) <= "00000000";
    MEMORY(097) <= "00000000";
    MEMORY(098) <= "00000000";
    MEMORY(099) <= "00000000";

    MEMORY(100) <= "00000000";
    MEMORY(101) <= "00000000";
    MEMORY(102) <= "00000000";
    MEMORY(103) <= "00000000";

    MEMORY(104) <= "00000000";
    MEMORY(105) <= "00000000";
    MEMORY(106) <= "00000000";
    MEMORY(107) <= "00000000";

    MEMORY(108) <= "00000000";
    MEMORY(109) <= "00000000";
    MEMORY(110) <= "00000000";
    MEMORY(111) <= "00000000";

    MEMORY(112) <= "00000000";
    MEMORY(113) <= "00000000";
    MEMORY(114) <= "00000000";
    MEMORY(115) <= "00000000";

    MEMORY(116) <= "00000000";
    MEMORY(117) <= "00000000";
    MEMORY(118) <= "00000000";
    MEMORY(119) <= "00000000";

    MEMORY(120) <= "00000000";
    MEMORY(121) <= "00000000";
    MEMORY(122) <= "00000000";
    MEMORY(123) <= "00000000";

    MEMORY(124) <= "00000000";
    MEMORY(125) <= "00000000";
    MEMORY(126) <= "00000000";
    MEMORY(127) <= "00000000";

    MEMORY(128) <= "00000000";
    MEMORY(129) <= "00000000";
    MEMORY(130) <= "00000000";
    MEMORY(131) <= "00000000";

    MEMORY(132) <= "00000000";
    MEMORY(133) <= "00000000";
    MEMORY(134) <= "00000000";
    MEMORY(135) <= "00000000";

    MEMORY(136) <= "00000000";
    MEMORY(137) <= "00000000";
    MEMORY(138) <= "00000000";
    MEMORY(139) <= "00000000";

    MEMORY(141) <= "00000000";
    MEMORY(142) <= "00000000";
    MEMORY(143) <= "00000000";
    MEMORY(144) <= "00000000";

    MEMORY(145) <= "00000000";
    MEMORY(146) <= "00000000";
    MEMORY(147) <= "00000000";
    MEMORY(148) <= "00000000";

    MEMORY(149) <= "00000000";
    MEMORY(150) <= "00000000";
    MEMORY(151) <= "00000000";
    MEMORY(152) <= "00000000";

    MEMORY(153) <= "00000000";
    MEMORY(154) <= "00000000";
    MEMORY(155) <= "00000000";
    MEMORY(156) <= "00000000";

    MEMORY(157) <= "00000000";
    MEMORY(158) <= "00000000";
    MEMORY(159) <= "00000000";
    MEMORY(160) <= "00000000";

    MEMORY(161) <= "00000000";
    MEMORY(162) <= "00000000";
    MEMORY(163) <= "00000000";
    MEMORY(164) <= "00000000";

    MEMORY(165) <= "00000000";
    MEMORY(166) <= "00000000";
    MEMORY(167) <= "00000000";
    MEMORY(168) <= "00000000";

    MEMORY(169) <= "00000000";
    MEMORY(170) <= "00000000";
    MEMORY(171) <= "00000000";
    MEMORY(172) <= "00000000";

    MEMORY(173) <= "00000000";
    MEMORY(174) <= "00000000";
    MEMORY(175) <= "00000000";
    MEMORY(176) <= "00000000";

    MEMORY(177) <= "00000000";
    MEMORY(178) <= "00000000";
    MEMORY(179) <= "00000000";
    MEMORY(180) <= "00000000";

    MEMORY(181) <= "00000000";
    MEMORY(182) <= "00000000";
    MEMORY(183) <= "00000000";
    MEMORY(184) <= "00000000";

    MEMORY(185) <= "00000000";
    MEMORY(186) <= "00000000";
    MEMORY(187) <= "00000000";
    MEMORY(188) <= "00000000";

    MEMORY(189) <= "00000000";
    MEMORY(190) <= "00000000";
    MEMORY(191) <= "00000000";
    MEMORY(192) <= "00000000";

    MEMORY(193) <= "00000000";
    MEMORY(194) <= "00000000";
    MEMORY(195) <= "00000000";
    MEMORY(196) <= "00000000";

    MEMORY(197) <= "00000000";
    MEMORY(198) <= "00000000";
    MEMORY(199) <= "00000000";
    MEMORY(200) <= "00000000";

    MEMORY(201) <= "00000000";
    MEMORY(202) <= "00000000";
    MEMORY(203) <= "00000000";
    MEMORY(204) <= "00000000";

    MEMORY(205) <= "00000000";
    MEMORY(206) <= "00000000";
    MEMORY(207) <= "00000000";
    MEMORY(208) <= "00000000";

    MEMORY(209) <= "00000000";
    MEMORY(210) <= "00000000";
    MEMORY(211) <= "00000000";
    MEMORY(212) <= "00000000";

    MEMORY(213) <= "00000000";
    MEMORY(214) <= "00000000";
    MEMORY(215) <= "00000000";
    MEMORY(216) <= "00000000";

    MEMORY(217) <= "00000000";
    MEMORY(218) <= "00000000";
    MEMORY(219) <= "00000000";
    MEMORY(220) <= "00000000";

    MEMORY(221) <= "00000000";
    MEMORY(222) <= "00000000";
    MEMORY(223) <= "00000000";
    MEMORY(224) <= "00000000";

    MEMORY(225) <= "00000000";
    MEMORY(226) <= "00000000";
    MEMORY(227) <= "00000000";
    MEMORY(228) <= "00000000";

    MEMORY(229) <= "00000000";
    MEMORY(230) <= "00000000";
    MEMORY(231) <= "00000000";
    MEMORY(232) <= "00000000";

    MEMORY(233) <= "00000000";
    MEMORY(234) <= "00000000";
    MEMORY(235) <= "00000000";
    MEMORY(236) <= "00000000";

    MEMORY(237) <= "00000000";
    MEMORY(238) <= "00000000";
    MEMORY(239) <= "00000000";
    MEMORY(240) <= "00000000";

    MEMORY(241) <= "00000000";
    MEMORY(242) <= "00000000";
    MEMORY(243) <= "00000000";
    MEMORY(244) <= "00000000";

    MEMORY(245) <= "00000000";
    MEMORY(246) <= "00000000";
    MEMORY(247) <= "00000000";
    MEMORY(248) <= "00000000";

    MEMORY(249) <= "00000000";
    MEMORY(250) <= "00000000";
    MEMORY(251) <= "00000000";
    MEMORY(252) <= "00000000";

    MEMORY(253) <= "00000000";
    MEMORY(254) <= "00000000";
    MEMORY(255) <= "00000000";
    MEMORY(256) <= "00000000";

    MEMORY(257) <= "00000000";
    MEMORY(258) <= "00000000";
    MEMORY(259) <= "00000000";
    MEMORY(260) <= "00000000";

    MEMORY(261) <= "00000000";
    MEMORY(262) <= "00000000";
    MEMORY(263) <= "00000000";
    MEMORY(264) <= "00000000";

    MEMORY(265) <= "00000000";
    MEMORY(266) <= "00000000";
    MEMORY(267) <= "00000000";
    MEMORY(268) <= "00000000";

    MEMORY(269) <= "00000000";
    MEMORY(270) <= "00000000";
    MEMORY(271) <= "00000000";
    MEMORY(272) <= "00000000";

    MEMORY(273) <= "00000000";
    MEMORY(274) <= "00000000";
    MEMORY(275) <= "00000000";
    MEMORY(276) <= "00000000";

    MEMORY(277) <= "00000000";
    MEMORY(278) <= "00000000";
    MEMORY(279) <= "00000000";
    MEMORY(280) <= "00000000";

    MEMORY(281) <= "00000000";
    MEMORY(282) <= "00000000";
    MEMORY(283) <= "00000000";
    MEMORY(284) <= "00000000";

    MEMORY(285) <= "00000000";
    MEMORY(286) <= "00000000";
    MEMORY(287) <= "00000000";
    MEMORY(288) <= "00000000";

    MEMORY(289) <= "00000000";
    MEMORY(290) <= "00000000";
    MEMORY(291) <= "00000000";
    MEMORY(292) <= "00000000";

    MEMORY(293) <= "00000000";
    MEMORY(294) <= "00000000";
    MEMORY(295) <= "00000000";
    MEMORY(296) <= "00000000";

    MEMORY(297) <= "00000000";
    MEMORY(298) <= "00000000";
    MEMORY(299) <= "00000000";
    MEMORY(300) <= "00000000";

    MEMORY(301) <= "00000000";
    MEMORY(302) <= "00000000";
    MEMORY(303) <= "00000000";
    MEMORY(304) <= "00000000";

    MEMORY(305) <= "00000000";
    MEMORY(306) <= "00000000";
    MEMORY(307) <= "00000000";
    MEMORY(308) <= "00000000";

    MEMORY(309) <= "00000000";
    MEMORY(310) <= "00000000";
    MEMORY(311) <= "00000000";
    MEMORY(312) <= "00000000";

    MEMORY(313) <= "00000000";
    MEMORY(314) <= "00000000";
    MEMORY(315) <= "00000000";
    MEMORY(316) <= "00000000";

    MEMORY(317) <= "00000000";
    MEMORY(318) <= "00000000";
    MEMORY(319) <= "00000000";
    MEMORY(320) <= "00000000";

    MEMORY(321) <= "00000000";
    MEMORY(322) <= "00000000";
    MEMORY(323) <= "00000000";
    MEMORY(324) <= "00000000";

    MEMORY(325) <= "00000000";
    MEMORY(326) <= "00000000";
    MEMORY(327) <= "00000000";
    MEMORY(328) <= "00000000";

    MEMORY(329) <= "00000000";
    MEMORY(330) <= "00000000";
    MEMORY(331) <= "00000000";
    MEMORY(332) <= "00000000";

    MEMORY(333) <= "00000000";
    MEMORY(334) <= "00000000";
    MEMORY(335) <= "00000000";
    MEMORY(336) <= "00000000";

    MEMORY(337) <= "00000000";
    MEMORY(338) <= "00000000";
    MEMORY(339) <= "00000000";
    MEMORY(340) <= "00000000";

    MEMORY(341) <= "00000000";
    MEMORY(342) <= "00000000";
    MEMORY(343) <= "00000000";
    MEMORY(344) <= "00000000";

    MEMORY(345) <= "00000000";
    MEMORY(346) <= "00000000";
    MEMORY(347) <= "00000000";
    MEMORY(348) <= "00000000";

    MEMORY(349) <= "00000000";
    MEMORY(350) <= "00000000";
    MEMORY(351) <= "00000000";
    MEMORY(352) <= "00000000";

    MEMORY(353) <= "00000000";
    MEMORY(354) <= "00000000";
    MEMORY(355) <= "00000000";
    MEMORY(356) <= "00000000";

    MEMORY(357) <= "00000000";
    MEMORY(358) <= "00000000";
    MEMORY(359) <= "00000000";
    MEMORY(360) <= "00000000";

    MEMORY(361) <= "00000000";
    MEMORY(362) <= "00000000";
    MEMORY(363) <= "00000000";
    MEMORY(364) <= "00000000";

    MEMORY(365) <= "00000000";
    MEMORY(366) <= "00000000";
    MEMORY(367) <= "00000000";
    MEMORY(368) <= "00000000";

    MEMORY(369) <= "00000000";
    MEMORY(370) <= "00000000";
    MEMORY(371) <= "00000000";
    MEMORY(372) <= "00000000";

    MEMORY(373) <= "00000000";
    MEMORY(374) <= "00000000";
    MEMORY(375) <= "00000000";
    MEMORY(376) <= "00000000";

    MEMORY(377) <= "00000000";
    MEMORY(378) <= "00000000";
    MEMORY(379) <= "00000000";
    MEMORY(380) <= "00000000";

    MEMORY(381) <= "00000000";
    MEMORY(382) <= "00000000";
    MEMORY(383) <= "00000000";
    MEMORY(384) <= "00000000";

    MEMORY(385) <= "00000000";
    MEMORY(386) <= "00000000";
    MEMORY(387) <= "00000000";
    MEMORY(388) <= "00000000";

    MEMORY(389) <= "00000000";
    MEMORY(390) <= "00000000";
    MEMORY(391) <= "00000000";
    MEMORY(392) <= "00000000";

    MEMORY(393) <= "00000000";
    MEMORY(394) <= "00000000";
    MEMORY(395) <= "00000000";
    MEMORY(396) <= "00000000";

    MEMORY(397) <= "00000000";
    MEMORY(398) <= "00000000";
    MEMORY(399) <= "00000000";
    MEMORY(400) <= "00000000";

    PROCESS (ADDRESS)
    BEGIN
        INSTRUCTION <=  MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))    ) &
                        MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1) &
                        MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 2) &
                        MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 3);
    END PROCESS;
END;