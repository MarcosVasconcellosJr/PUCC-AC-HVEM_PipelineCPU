LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Cpu IS
    GENERIC (DATA_SIZE : INTEGER := 32); -- Generic data size to map in components
    PORT (
        CLOCK : IN STD_LOGIC;
        INSTRUCTION_OUT_IFID : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_REGS_PC : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_CONTROL : OUT STD_LOGIC;
        DEB_ULA_IN_1 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_ULA_IN_2 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_OUT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_RegDst : OUT STD_LOGIC_VECTOR(0 TO 4);

        DEB_REG_ULA_IN_1 : OUT STD_LOGIC_VECTOR(0 TO 4);

        DEB_SINAL_MUX_MEMWB : OUT STD_LOGIC;
        DEB_SINAL_REG_WRITE : OUT STD_LOGIC;
        DEB_WRITE_REG : OUT STD_LOGIC_VECTOR(0 TO 4);
        DEB_WRITE_DATA : OUT STD_LOGIC_VECTOR(0 TO 31);

        DEB_FILE_REG_1 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_FILE_REG_2 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_FILE_REG_3 : OUT STD_LOGIC_VECTOR(0 TO 31);
        DEB_FILE_REG_AUX : OUT STD_LOGIC
    );
END Cpu;
ARCHITECTURE CPU OF Cpu IS

    -- ControlUnit - PORT MAP
    COMPONENT ControlUnit
        PORT (
            WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            EX : OUT STD_LOGIC_VECTOR(0 TO 4);
            SIGNAL_JUMP : OUT STD_LOGIC_VECTOR(0 TO 1);
            INSTRUCTION : IN STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- AluControl - PORT MAP
    COMPONENT AluControl
        PORT (
            ALU_OP : IN STD_LOGIC_VECTOR(0 TO 2);
            FUNCT : IN STD_LOGIC_VECTOR(0 TO 5);
            ULA_CODE : OUT STD_LOGIC_VECTOR(0 TO 1)
        );
    END COMPONENT;

    -- ShiftLeft - PORT MAP
    COMPONENT ShiftLeft
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 31);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- ShiftLeft2_26to28 - PORT MAP
    COMPONENT ShiftLeft2_26to28
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 25);
            X : OUT STD_LOGIC_VECTOR(0 TO 27)
        );
    END COMPONENT;

    -- Signal Extend - PORT MAP
    COMPONENT SignalExtend
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 15);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- Mux_2to1_32b - PORT MAP
    COMPONENT Mux_2to1_32b
        PORT (
            CONTROL : IN STD_LOGIC;
            A : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
            B : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);
            X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1)
        );
    END COMPONENT;

    --  Generic3to1Mux - PORT MAP
    COMPONENT Generic3to1Mux
        PORT (
            JUMP_SIGNAL : IN STD_LOGIC_VECTOR (0 TO 1);
            A, B, C : IN STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1);

            X : OUT STD_LOGIC_VECTOR (0 TO DATA_SIZE - 1)
        );
    END COMPONENT;

    -- Alu - PORT MAP
    COMPONENT Alu
        PORT (
            A : IN STD_LOGIC_VECTOR(0 TO 31);
            B : IN STD_LOGIC_VECTOR(0 TO 31);
            ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1);
            ALU_OUT : OUT STD_LOGIC_VECTOR(0 TO 31);
            ZERO : OUT STD_LOGIC
        );
    END COMPONENT;

    -- Data Memory - PORT MAP
    COMPONENT DataMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
            CLOCK : IN STD_LOGIC;
            MEM_WRITE : IN STD_LOGIC;
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 31);
            MEM_READ : IN STD_LOGIC;
            READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- InstructionMemory - PORT MAP
    COMPONENT InstructionMemory
        PORT (
            ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
            INSTRUCTION : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"
        );
    END COMPONENT;

    -- PCIncrement - PORT MAP
    COMPONENT PCIncrement
        PORT (
            PC : IN STD_LOGIC_VECTOR (0 TO 31);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- Reg_Pipe_IFID - PORT MAP
    COMPONENT Reg_Pipe_IFID
        PORT (
            CLOCK : IN STD_LOGIC;
            IN_PC_MAIS_4 : IN STD_LOGIC_VECTOR(0 TO 31);
            IN_INSTR_MEM : IN STD_LOGIC_VECTOR(0 TO 31);

            OUT_PC_MAIS_4 : OUT STD_LOGIC_VECTOR(0 TO 31);
            OUT_INSTR_MEM : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- Mux_2to1_5b - PORT MAP
    COMPONENT Mux_2to1_5b
        PORT (
            CONTROL : IN STD_LOGIC; -- Controller to select the desired data
            A : IN STD_LOGIC_VECTOR (0 TO 4); -- The first data option
            B : IN STD_LOGIC_VECTOR (0 TO 4); -- The second data option
            X : OUT STD_LOGIC_VECTOR (0 TO 4)
        );

    END COMPONENT;

    -- Reg_Pipe_IDEX - PORT MAP
    COMPONENT Reg_Pipe_IDEX
        PORT (
            CLOCK : IN STD_LOGIC;
            IDEX_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            IDEX_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            IDEX_IN_EX : IN STD_LOGIC_VECTOR(0 TO 4);
            IDEX_IN_PC : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_READ1 : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_IMED : IN STD_LOGIC_VECTOR(0 TO 31);
            IDEX_IN_RT : IN STD_LOGIC_VECTOR(0 TO 4);
            IDEX_IN_RD : IN STD_LOGIC_VECTOR(0 TO 4);

            IDEX_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            IDEX_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            IDEX_OUT_EX : OUT STD_LOGIC_VECTOR(0 TO 4);
            IDEX_OUT_PC : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_READ1 : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_IMED : OUT STD_LOGIC_VECTOR(0 TO 31);
            IDEX_OUT_RT : OUT STD_LOGIC_VECTOR(0 TO 4);
            IDEX_OUT_RD : OUT STD_LOGIC_VECTOR(0 TO 4)
        );
    END COMPONENT;

    -- Reg_Pipe_EXMEM - PORT MAP
    COMPONENT Reg_Pipe_EXMEM
        PORT (
            CLOCK : IN STD_LOGIC;
            EXMEM_IN_ZERO : IN STD_LOGIC;
            EXMEM_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_IN_MEM : IN STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_IN_RESULT_ADDER : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_READ2 : IN STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 4);

            EXMEM_OUT_ZERO : OUT STD_LOGIC;
            EXMEM_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            EXMEM_OUT_MEM : OUT STD_LOGIC_VECTOR(0 TO 2);
            EXMEM_OUT_RESULT_ADDER : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_READ2 : OUT STD_LOGIC_VECTOR(0 TO 31);
            EXMEM_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 4)
        );
    END COMPONENT;

    -- Reg_Pipe_MEMWB - PORT MAP
    COMPONENT Reg_Pipe_MEMWB
        PORT (
            CLOCK : IN STD_LOGIC;
            MEMWB_IN_WB : IN STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_IN_RESULT_ULA : IN STD_LOGIC_VECTOR(0 TO 31);
            MEMWB_IN_REGDST : IN STD_LOGIC_VECTOR(0 TO 4);
            MEMWB_IN_READ_DATA : IN STD_LOGIC_VECTOR(0 TO 31);

            MEMWB_OUT_WB : OUT STD_LOGIC_VECTOR(0 TO 1);
            MEMWB_OUT_RESULT_ULA : OUT STD_LOGIC_VECTOR(0 TO 31);
            MEMWB_OUT_REGDST : OUT STD_LOGIC_VECTOR(0 TO 4);
            MEMWB_OUT_READ_DATA : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- FileRegister - PORT MAP
    COMPONENT FileRegister
        PORT (
            REGWRITE : IN STD_LOGIC;
            CLOCK : IN STD_LOGIC;
            READ_REGISTER_1 : IN STD_LOGIC_VECTOR(0 TO 4);
            READ_REGISTER_2 : IN STD_LOGIC_VECTOR(0 TO 4);
            WRITE_REGISTER : IN STD_LOGIC_VECTOR(0 TO 4);
            WRITE_DATA : IN STD_LOGIC_VECTOR(0 TO 31);

            READ_DATA_1 : OUT STD_LOGIC_VECTOR(0 TO 31);
            READ_DATA_2 : OUT STD_LOGIC_VECTOR(0 TO 31);

            DEB_FILE_REG_1 : OUT STD_LOGIC_VECTOR(0 TO 31);

            DEB_FILE_REG_2 : OUT STD_LOGIC_VECTOR(0 TO 31);
            DEB_FILE_REG_3 : OUT STD_LOGIC_VECTOR(0 TO 31);
            DEB_FILE_REG_AUX : OUT STD_LOGIC
        );
    END COMPONENT;

    -- FileRegister - PORT MAP
    COMPONENT ProgramCounter
        PORT (
            CLOCK : IN STD_LOGIC;
            PC_INC : IN STD_LOGIC_VECTOR(0 TO 31);
            PC : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    -- SignExtend - PORT MAP
    COMPONENT SignExtend
        PORT (
            A : IN STD_LOGIC_VECTOR (0 TO 15);
            X : OUT STD_LOGIC_VECTOR(0 TO 31)
        );
    END COMPONENT;

    ---------------------------------------------------------------------------------------------------------------
    --------------------------------------------------- SIGNALS ---------------------------------------------------

    -- Used to do nothing normally
    SIGNAL UNUSED : STD_LOGIC;

    --******************** INSTRUCTION FETCH ********************--

    -- SIGNALS - TO CONTROL COMPONENT INTERACTION IN EXECUTION TIME
    SIGNAL SIG_PC_SRC : STD_LOGIC;
    SIGNAL SIG_JUMP : STD_LOGIC;

    -- WIRES - TO CONNECT PORT MAP BETWEEN COMPONENTS
    SIGNAL WIRE_OUT_PC_INC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_PC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_PC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_JUMP : STD_LOGIC_VECTOR(0 TO 31); --Used to connect mux 
    SIGNAL WIRE_INST_MEM_IFID : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_PC_PC : STD_LOGIC_VECTOR(0 TO 31);

    SIGNAL WIRE_SHIFT_MUX_JUMP : STD_LOGIC_VECTOR(0 TO 27);
    SIGNAL WIRE_SHIFT_CONCAT : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_PC_MUX_JUMP : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_JUMP_PC : STD_LOGIC_VECTOR(0 TO 31);
    ---------------------------------------------------------------------------------------------------------------
    --------------------------------------------------- DECODE STAGE ---------------------------------------------------

    --WIRES
    SIGNAL WIRE_PC_INC_IFID_TO_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_IFID_INSTRUCTION : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_READ_DATA1_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_READ_DATA2_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_SIGNAL_EXTEND_IDEX : STD_LOGIC_VECTOR(0 TO 31);
    -- Control Unit
    SIGNAL WIRE_UC_IDEX_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_UC_IDEX_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_UC_IDEX_EX : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_UC_JUMP_SIGNAL : STD_LOGIC_VECTOR(0 TO 1) := "00";

    --******************** INSTRUCTION EXECUTION STAGE  ********************--

    -- WIRES OF REG_PIPE
    SIGNAL WIRE_IDEX_WB_EXMEM_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_IDEX_MEM_EXMEM_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_PC_INC_IDEX_TO_ADDER : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_READ1_ALU_A : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_IDEX_READ2 : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_IDEX_IMED : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_IDEX_RT_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_IDEX_RD_MUX_REGDST : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_OUT_IDEX_EX : STD_LOGIC_VECTOR(0 TO 4);
    -- WIRES OF THIS STAGE
    SIGNAL WIRE_SHIFT_LEFT_ADDER_B : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_ALU_B : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MUX_REGDST_EXMEM : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_ULA_CODE : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_ALU_RES_EXMEM : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_ZERO_EXMEM : STD_LOGIC;
    SIGNAL WIRE_ADDER_RES_EXMEM : STD_LOGIC_VECTOR(0 TO 31);

    --******************** INSTRUCTION MEMORY STAGE ********************--

    -- WIRES OF REG_PIPE
    SIGNAL WIRE_OUT_EXMEM_ZERO : STD_LOGIC;
    SIGNAL WIRE_EXMEM_WB_MEMWB_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_OUT_EXMEM_MEM : STD_LOGIC_VECTOR(0 TO 2);
    SIGNAL WIRE_EXMEM_ADDER_RES_MUXPC : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_OUT_EXMEM_ALU_RES : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_EXMEM_READ2_WRITE_DATA : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_EXMEM_REGDST_MEM_WB : STD_LOGIC_VECTOR(0 TO 4);

    -- WIRES OF THIS STAGE

    SIGNAL PCSrc : STD_LOGIC := '0';
    SIGNAL WIRE_READ_DATA_MEMWB : STD_LOGIC_VECTOR(0 TO 31);

    --******************** INSTRUCTION WRITE BACK STAGE ********************--

    -- WIRES OF REG_PIPE
    SIGNAL WIRE_OUT_MEMWB_WB : STD_LOGIC_VECTOR(0 TO 1);
    SIGNAL WIRE_MEMWB_ALU_RES : STD_LOGIC_VECTOR(0 TO 31);
    SIGNAL WIRE_MEMWB_REG_DST : STD_LOGIC_VECTOR(0 TO 4);
    SIGNAL WIRE_MEMWB_READ_DATA_MUX_WB : STD_LOGIC_VECTOR(0 TO 31);
    --
    SIGNAL WIRE_MUX_WB_WRITE_DATA : STD_LOGIC_VECTOR(0 TO 31);

BEGIN

    --******************** COMPONENTS INSTRUCTION FETCH ********************--

    INST_MEM : InstructionMemory PORT MAP(WIRE_OUT_PC, WIRE_INST_MEM_IFID);
    MUX_PC : Mux_2to1_32b PORT MAP(PCSrc, WIRE_OUT_PC_INC, WIRE_EXMEM_ADDER_RES_MUXPC, WIRE_MUX_PC_MUX_JUMP);
    PC_INC : PCIncrement PORT MAP(WIRE_OUT_PC, WIRE_OUT_PC_INC);
    MUX_JUMP : Generic3to1Mux PORT MAP(WIRE_UC_JUMP_SIGNAL, WIRE_MUX_PC_MUX_JUMP, WIRE_SHIFT_CONCAT, WIRE_READ_DATA1_IDEX, WIRE_MUX_JUMP_PC);
    PC : ProgramCounter PORT MAP(CLOCK, WIRE_MUX_JUMP_PC, WIRE_OUT_PC);

    DEB_REGS_PC <= WIRE_OUT_PC_INC;
    --******************** REG_PIPELINE IF/ID ********************--

    IFID : Reg_Pipe_IFID PORT MAP(CLOCK, WIRE_OUT_PC_INC, WIRE_INST_MEM_IFID, WIRE_PC_INC_IFID_TO_IDEX, WIRE_OUT_IFID_INSTRUCTION);

    INSTRUCTION_OUT_IFID <= WIRE_OUT_IFID_INSTRUCTION;

    --******************** COMPONENTS INSTRUCTION DECODE STAGE ********************--

    WIRE_SHIFT_CONCAT <= WIRE_SHIFT_MUX_JUMP & WIRE_PC_INC_IFID_TO_IDEX(0 TO 3);

    SHIFT_IF : ShiftLeft2_26to28 PORT MAP(WIRE_OUT_IFID_INSTRUCTION(0 TO 25), WIRE_SHIFT_MUX_JUMP);

    DEB_REG_ULA_IN_1 <= WIRE_OUT_IFID_INSTRUCTION(6 TO 10);
    DEB_SINAL_REG_WRITE <= WIRE_OUT_MEMWB_WB(0);
    FILE_REG : FileRegister PORT MAP(
        WIRE_OUT_MEMWB_WB(0),
        CLOCK,
        WIRE_OUT_IFID_INSTRUCTION(6 TO 10),
        WIRE_OUT_IFID_INSTRUCTION(11 TO 15),
        WIRE_MEMWB_REG_DST,
        WIRE_MUX_WB_WRITE_DATA,
        WIRE_READ_DATA1_IDEX,
        WIRE_READ_DATA2_IDEX,

        DEB_FILE_REG_1,
        DEB_FILE_REG_2,
        DEB_FILE_REG_3,

        DEB_FILE_REG_AUX
    );
    SIGNAL_EXTEND : SignExtend PORT MAP(WIRE_OUT_IFID_INSTRUCTION(16 TO 31), WIRE_SIGNAL_EXTEND_IDEX);
    UC : ControlUnit PORT MAP(WIRE_UC_IDEX_WB, WIRE_UC_IDEX_MEM, WIRE_UC_IDEX_EX, WIRE_UC_JUMP_SIGNAL, WIRE_OUT_IFID_INSTRUCTION);

    --******************** REG_PIPELINE ID/EX ********************--
    IDEX : Reg_Pipe_IDEX PORT MAP(
        -- IN --
        CLOCK, WIRE_UC_IDEX_WB, WIRE_UC_IDEX_MEM, WIRE_UC_IDEX_EX, WIRE_PC_INC_IFID_TO_IDEX, WIRE_READ_DATA1_IDEX, WIRE_READ_DATA2_IDEX, WIRE_SIGNAL_EXTEND_IDEX, WIRE_OUT_IFID_INSTRUCTION(11 TO 15), WIRE_OUT_IFID_INSTRUCTION(16 TO 20),
        -- OUT --
        WIRE_IDEX_WB_EXMEM_WB, WIRE_IDEX_MEM_EXMEM_MEM, WIRE_OUT_IDEX_EX, WIRE_PC_INC_IDEX_TO_ADDER, WIRE_IDEX_READ1_ALU_A, WIRE_OUT_IDEX_READ2, WIRE_OUT_IDEX_IMED, WIRE_IDEX_RT_MUX_REGDST, WIRE_IDEX_RD_MUX_REGDST
    );
    --******************** COMPONENTS INSTRUCTION EXECUTION  ********************--

    SHIFT_LEFT : ShiftLeft PORT MAP(WIRE_OUT_IDEX_IMED, WIRE_SHIFT_LEFT_ADDER_B);
    MUX_ALU_B : Mux_2to1_32b PORT MAP(WIRE_OUT_IDEX_EX(4), WIRE_OUT_IDEX_READ2, WIRE_OUT_IDEX_IMED, WIRE_MUX_ALU_B);
    MUX_REGDST : Mux_2to1_5b PORT MAP(WIRE_OUT_IDEX_EX(0), WIRE_IDEX_RT_MUX_REGDST, WIRE_IDEX_RD_MUX_REGDST, WIRE_MUX_REGDST_EXMEM);
    ALU_CONTROL : AluControl PORT MAP(WIRE_OUT_IDEX_EX(1 TO 3), WIRE_OUT_IDEX_IMED(26 TO 31), WIRE_ULA_CODE);
    ADDER_SHIFT2_PC_INC : Alu PORT MAP(WIRE_PC_INC_IDEX_TO_ADDER, WIRE_SHIFT_LEFT_ADDER_B, "00", WIRE_ADDER_RES_EXMEM, UNUSED);
    MAIN_ALU : Alu PORT MAP(WIRE_IDEX_READ1_ALU_A, WIRE_MUX_ALU_B, WIRE_ULA_CODE, WIRE_ALU_RES_EXMEM, WIRE_ZERO_EXMEM);

    DEB_CONTROL <= WIRE_OUT_IDEX_EX(0);
    DEB_ULA_IN_1 <= WIRE_IDEX_READ1_ALU_A;
    DEB_ULA_IN_2 <= WIRE_MUX_ALU_B;
    DEB_OUT_ULA <= WIRE_ALU_RES_EXMEM;
    DEB_RegDst <= WIRE_MUX_REGDST_EXMEM;
    --******************** REG_PIPELINE EX/MEM ********************--
    EXMEM : Reg_Pipe_EXMEM PORT MAP(
        -- IN --
        CLOCK,
        WIRE_ZERO_EXMEM,
        WIRE_IDEX_WB_EXMEM_WB,
        WIRE_IDEX_MEM_EXMEM_MEM,
        WIRE_ADDER_RES_EXMEM,
        WIRE_ALU_RES_EXMEM,
        WIRE_OUT_IDEX_READ2,
        WIRE_MUX_REGDST_EXMEM,
        -- OUT --
        WIRE_OUT_EXMEM_ZERO,
        WIRE_EXMEM_WB_MEMWB_WB,
        WIRE_OUT_EXMEM_MEM,
        WIRE_EXMEM_ADDER_RES_MUXPC,
        WIRE_OUT_EXMEM_ALU_RES,
        WIRE_EXMEM_READ2_WRITE_DATA,
        WIRE_EXMEM_REGDST_MEM_WB
    );

    --******************** COMPONENTS INSTRUCTION MEMORY  ********************--
    PCSrc <= WIRE_OUT_EXMEM_MEM(0) AND WIRE_OUT_EXMEM_ZERO;
    DATA_MEMORY : DataMemory PORT MAP(WIRE_OUT_EXMEM_ALU_RES, CLOCK, WIRE_OUT_EXMEM_MEM(2), WIRE_EXMEM_READ2_WRITE_DATA, WIRE_OUT_EXMEM_MEM(1), WIRE_READ_DATA_MEMWB);

    --******************** REG_PIPELINE MEM/WB ********************--

    MEMWB : Reg_Pipe_MEMWB PORT MAP(
        -- IN --
        CLOCK,
        WIRE_EXMEM_WB_MEMWB_WB,
        WIRE_OUT_EXMEM_ALU_RES,
        WIRE_EXMEM_REGDST_MEM_WB,
        WIRE_READ_DATA_MEMWB,
        -- OUT --
        WIRE_OUT_MEMWB_WB,
        WIRE_MEMWB_ALU_RES,
        WIRE_MEMWB_REG_DST,
        WIRE_MEMWB_READ_DATA_MUX_WB
    );

    --******************** COMPONENTS INSTRUCTION WRITE BACK ********************--
    MUX_WB : Mux_2to1_32b PORT MAP(WIRE_OUT_MEMWB_WB(1), WIRE_MEMWB_READ_DATA_MUX_WB, WIRE_MEMWB_ALU_RES, WIRE_MUX_WB_WRITE_DATA);
    DEB_SINAL_MUX_MEMWB <= WIRE_OUT_MEMWB_WB(1);

    DEB_WRITE_REG <= WIRE_MEMWB_REG_DST;
    DEB_WRITE_DATA <= WIRE_MUX_WB_WRITE_DATA;

    ---------------------------------------------------------------------------------------------------------------
    ---------------------------------------------------- DEBUG ----------------------------------------------------
END;