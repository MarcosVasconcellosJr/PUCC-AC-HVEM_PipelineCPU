LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Alu IS
	PORT (
		A : IN STD_LOGIC_VECTOR(0 TO 31); -- REGISTER
		B : IN STD_LOGIC_VECTOR(0 TO 31); -- REGISTER
		ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1); -- CODE OF THE ARITHMETIC OPERATION OPTION
		ALU_OUT : OUT STD_LOGIC_VECTOR(0 TO 31); -- WHERE WE WILL STORE THE RESULT OF THE ARITHMETIC OPERATION
		ZERO : OUT STD_LOGIC);
END Alu;

ARCHITECTURE ALU OF Alu IS
	SIGNAL AUX : STD_LOGIC_VECTOR(0 TO 31);
BEGIN
	PROCESS (A, B, ALU_CODE)
	BEGIN
		-- SWITCH CASE TO DO THE RIGHT OPERATION BASED IN ALU_CODE
		CASE ALU_CODE IS
			WHEN "00" => AUX <= A + B;
			WHEN "01" => AUX <= A - B;
			WHEN "10" => AUX <= A AND B;
			WHEN "11" => AUX <= A OR B;
			WHEN OTHERS => AUX <= "00000000000000000000000000000000";
		END CASE;
		IF (AUX = "00000000000000000000000000000000") THEN
			ZERO <= '1';
		ELSE
			ZERO <= '0';
		END IF;

		ALU_OUT <= AUX;
	END PROCESS;
END ALU;