LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ALU IS
	PORT (
		RS_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- REGISTER
		RS_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0); -- REGISTER
		ALU_CODE : IN STD_LOGIC_VECTOR(0 TO 1); -- CODE OF THE ARITHMETIC OPERATION OPTION
		ALU_OUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)); -- WHERE WE WILL STORE THE RESULT OF THE ARITHMETIC OPERATION
END ALU;

ARCHITECTURE ALU OF ALU IS
BEGIN
	PROCESS (RS_DATA, RS_DATA, ALU_CODE)
	BEGIN
		-- SWITCH CASE TO DO THE RIGHT OPERATION BASED IN ALU_CODE
		CASE ALU_CODE IS
			WHEN "00" => ALU_OUT <= RS_DATA + RS_DATA;
			WHEN "01" => ALU_OUT <= RS_DATA - RS_DATA;
			WHEN "10" => ALU_OUT <= RS_DATA AND RS_DATA;
			WHEN "11" => ALU_OUT <= RS_DATA OR RS_DATA;
			WHEN OTHERS => ALU_OUT <= "00000000000000000000000000000000";
		END CASE;
	END PROCESS;
END ALU;