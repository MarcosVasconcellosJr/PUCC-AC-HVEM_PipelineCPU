LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Generic2to1Mux IS
    GENERIC (DATA_SIZE : INTEGER := 32);
    PORT (
        CONTROL : IN STD_LOGIC;
        A : IN STD_LOGIC_VECTOR (DATA_SIZE - 1 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR (DATA_SIZE - 1 DOWNTO 0);
        X : OUT STD_LOGIC_VECTOR (DATA_SIZE - 1 DOWNTO 0));
END Generic2to1Mux;

ARCHITECTURE MUX OF Generic2to1Mux IS
BEGIN
    X <= A WHEN (CONTROL == '1') ELSE B;
END;