LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY InstructionMemory IS

    PORT (
        ADDRESS : IN STD_LOGIC_VECTOR(0 TO 31);
        INSTRUCTION : OUT STD_LOGIC_VECTOR(0 TO 31) := "00000000000000000000000000000000"
    );

END InstructionMemory;

ARCHITECTURE MEM OF InstructionMemory IS
    TYPE MEM_TYPE IS ARRAY(0 TO 400) OF STD_LOGIC_VECTOR(0 TO 7);
    SIGNAL MEMORY : MEM_TYPE;
BEGIN
    -- LOADED WITH:

    -- ADDI $2, $2, 8
    -- SW $2, 0($4)
    -- LW $3, 0($4)
    -- ADDI $3, $6, 0
    -- JR $3

    -- Expected result: Infinite 8 times table in $2 register

    -- MEMORY(000) <= "00001000";
    -- MEMORY(001) <= "01000010";
    -- MEMORY(002) <= "00000000";
    -- MEMORY(003) <= "00001000";
    --
    -- MEMORY(004) <= "00000000";
    -- MEMORY(005) <= "00000000";
    -- MEMORY(006) <= "00000000";
    -- MEMORY(007) <= "00000000";
    --
    -- MEMORY(008) <= "00000000";
    -- MEMORY(009) <= "00000000";
    -- MEMORY(010) <= "00000000";
    -- MEMORY(011) <= "00000000";
    --
    -- MEMORY(012) <= "00000000";
    -- MEMORY(013) <= "00000000";
    -- MEMORY(014) <= "00000000";
    -- MEMORY(015) <= "00000000";
    -- MEMORY(016) <= "00011100";

    -- MEMORY(017) <= "10000010";
    -- MEMORY(018) <= "00000000";
    -- MEMORY(019) <= "00000000";
    --
    -- MEMORY(020) <= "00000000";
    -- MEMORY(021) <= "00000000";
    -- MEMORY(022) <= "00000000";
    -- MEMORY(023) <= "00000000";
    --
    -- MEMORY(024) <= "00000000";
    -- MEMORY(025) <= "00000000";
    -- MEMORY(026) <= "00000000";
    -- MEMORY(027) <= "00000000";
    --
    -- MEMORY(028) <= "00000000";
    -- MEMORY(029) <= "00000000";
    -- MEMORY(030) <= "00000000";
    -- MEMORY(031) <= "00000000";
    -- MEMORY(032) <= "00011000";

    -- MEMORY(033) <= "10000011";
    -- MEMORY(034) <= "00000000";
    -- MEMORY(035) <= "00000000";
    --
    -- MEMORY(036) <= "00000000";
    -- MEMORY(037) <= "00000000";
    -- MEMORY(038) <= "00000000";
    -- MEMORY(039) <= "00000000";
    --
    -- MEMORY(040) <= "00000000";
    -- MEMORY(041) <= "00000000";
    -- MEMORY(042) <= "00000000";
    -- MEMORY(043) <= "00000000";
    --
    -- MEMORY(044) <= "00000000";
    -- MEMORY(045) <= "00000000";
    -- MEMORY(046) <= "00000000";
    -- MEMORY(047) <= "00000000";
    --
    -- MEMORY(048) <= "00000000";
    -- MEMORY(049) <= "00000000";
    -- MEMORY(050) <= "00000000";
    -- MEMORY(051) <= "00000000";
    --
    -- MEMORY(052) <= "00000000";
    -- MEMORY(053) <= "00000000";
    -- MEMORY(054) <= "00000000";
    -- MEMORY(055) <= "00000000";
    --
    -- MEMORY(056) <= "00000000";
    -- MEMORY(057) <= "00000000";
    -- MEMORY(058) <= "00000000";
    -- MEMORY(059) <= "00000000";

    -- MEMORY(060) <= "00001000";
    -- MEMORY(061) <= "11000011";
    -- MEMORY(062) <= "00000000";
    -- MEMORY(063) <= "00000000";
    --
    -- MEMORY(064) <= "00000000";
    -- MEMORY(065) <= "00000000";
    -- MEMORY(066) <= "00000000";
    -- MEMORY(067) <= "00000000";
    --
    -- MEMORY(068) <= "00000000";
    -- MEMORY(069) <= "00000000";
    -- MEMORY(070) <= "00000000";
    -- MEMORY(071) <= "00000000";
    --
    -- MEMORY(072) <= "00000000";
    -- MEMORY(073) <= "00000000";
    -- MEMORY(074) <= "00000000";
    -- MEMORY(075) <= "00000000";
    --
    -- MEMORY(076) <= "00000000";
    -- MEMORY(077) <= "00000000";
    -- MEMORY(078) <= "00000000";
    -- MEMORY(079) <= "00000000";

    -- MEMORY(080) <= "00101000";
    -- MEMORY(081) <= "01100000";
    -- MEMORY(082) <= "00000000";
    -- MEMORY(083) <= "00000000";

    ---------------------------------------------------------------------------------------

    -- LOADED WITH:

    -- ORI $1, $1, 5
    -- ADDI $3, $3, 7
    -- J NEXT_INSTR
    -- SUBI $4, $1, 1
    -- NEXT_INSTR:
    -- AND $3, $3, $1

    -- Expected result: 5 in register 3 and 0 in register 2

    MEMORY(000) <= "00010100";
    MEMORY(001) <= "00100001";
    MEMORY(002) <= "00000000";
    MEMORY(003) <= "00000101";

    MEMORY(004) <= "00000000";
    MEMORY(005) <= "00000000";
    MEMORY(006) <= "00000000";
    MEMORY(007) <= "00000000";

    MEMORY(008) <= "00000000";
    MEMORY(009) <= "00000000";
    MEMORY(010) <= "00000000";
    MEMORY(011) <= "00000000";

    MEMORY(012) <= "00000000";
    MEMORY(013) <= "00000000";
    MEMORY(014) <= "00000000";
    MEMORY(015) <= "00000000";

    MEMORY(016) <= "00000000";
    MEMORY(017) <= "00000000";
    MEMORY(018) <= "00000000";
    MEMORY(019) <= "00000000";

    MEMORY(020) <= "00001000";
    MEMORY(021) <= "01100011";
    MEMORY(022) <= "00000000";
    MEMORY(023) <= "00000111";

    MEMORY(024) <= "00000000";
    MEMORY(025) <= "00000000";
    MEMORY(026) <= "00000000";
    MEMORY(027) <= "00000000";

    MEMORY(028) <= "00000000";
    MEMORY(029) <= "00000000";
    MEMORY(030) <= "00000000";
    MEMORY(031) <= "00000000";

    MEMORY(032) <= "00000000";
    MEMORY(033) <= "00000000";
    MEMORY(034) <= "00000000";
    MEMORY(035) <= "00000000";

    MEMORY(036) <= "00100100";
    MEMORY(037) <= "00000000";
    MEMORY(038) <= "00000000";
    MEMORY(039) <= "00010011";

    MEMORY(040) <= "00000000";
    MEMORY(041) <= "00000000";
    MEMORY(042) <= "00000000";
    MEMORY(043) <= "00000000";

    MEMORY(044) <= "00000000";
    MEMORY(045) <= "00000000";
    MEMORY(046) <= "00000000";
    MEMORY(047) <= "00000000";

    MEMORY(048) <= "00000000";
    MEMORY(049) <= "00000000";
    MEMORY(050) <= "00000000";
    MEMORY(051) <= "00000000";

    MEMORY(052) <= "00000000";
    MEMORY(053) <= "00000000";
    MEMORY(054) <= "00000000";
    MEMORY(055) <= "00000000";

    MEMORY(056) <= "00001100";
    MEMORY(057) <= "00100010";
    MEMORY(058) <= "00000000";
    MEMORY(059) <= "00000001";

    MEMORY(060) <= "00000000";
    MEMORY(061) <= "00000000";
    MEMORY(062) <= "00000000";
    MEMORY(063) <= "00000000";

    MEMORY(064) <= "00000000";
    MEMORY(065) <= "00000000";
    MEMORY(066) <= "00000000";
    MEMORY(067) <= "00000000";

    MEMORY(068) <= "00000000";
    MEMORY(069) <= "00000000";
    MEMORY(070) <= "00000000";
    MEMORY(071) <= "00000000";

    MEMORY(072) <= "00000000";
    MEMORY(073) <= "00000000";
    MEMORY(074) <= "00000000";
    MEMORY(075) <= "00000000";

    MEMORY(076) <= "00000000";
    MEMORY(077) <= "00000000";
    MEMORY(078) <= "00000000";
    MEMORY(079) <= "00000000";

    MEMORY(080) <= "00000100";
    MEMORY(081) <= "01100001";
    MEMORY(082) <= "00011000";
    MEMORY(083) <= "00100100";

    ---------------------------------------------------------------------------------------

    -- LOADED WITH:

    --     ADDI $1, $1, 5
    -- ADD $2, $2, $1
    -- LOOP:
    --     ADDI $1, $1, 5
    --     ADDI $3, $3, 1
    --     BEQ $3, $2, J_SUB
    --     J LOOP
    -- J_SUB:
    --     SUB $1, $3, $1

    -- Expected result: 25 in $1 register

    -- MEMORY(000) <= "00001000";
    -- MEMORY(001) <= "00100001";
    -- MEMORY(002) <= "00000000";
    -- MEMORY(003) <= "00000101";
    -- 
    -- MEMORY(004) <= "00000000";
    -- MEMORY(005) <= "00000000";
    -- MEMORY(006) <= "00000000";
    -- MEMORY(007) <= "00000000";
    -- 
    -- MEMORY(008) <= "00000000";
    -- MEMORY(009) <= "00000000";
    -- MEMORY(010) <= "00000000";
    -- MEMORY(011) <= "00000000";
    -- 
    -- MEMORY(012) <= "00000000";
    -- MEMORY(013) <= "00000000";
    -- MEMORY(014) <= "00000000";
    -- MEMORY(015) <= "00000000";
    -- 
    -- MEMORY(016) <= "00000100";
    -- MEMORY(017) <= "01000001";
    -- MEMORY(018) <= "00010000";
    -- MEMORY(019) <= "00100000";
    -- 
    -- MEMORY(020) <= "00000000";
    -- MEMORY(021) <= "00000000";
    -- MEMORY(022) <= "00000000";
    -- MEMORY(023) <= "00000000";
    -- 
    -- MEMORY(024) <= "00000000";
    -- MEMORY(025) <= "00000000";
    -- MEMORY(026) <= "00000000";
    -- MEMORY(027) <= "00000000";
    -- 
    -- MEMORY(028) <= "00000000";
    -- MEMORY(029) <= "00000000";
    -- MEMORY(030) <= "00000000";
    -- MEMORY(031) <= "00000000";
    -- 
    -- MEMORY(032) <= "00001000";
    -- MEMORY(033) <= "00100001";
    -- MEMORY(034) <= "00000000";
    -- MEMORY(035) <= "00000101";
    -- 
    -- MEMORY(036) <= "00000000";
    -- MEMORY(037) <= "00000000";
    -- MEMORY(038) <= "00000000";
    -- MEMORY(039) <= "00000000";
    -- 
    -- MEMORY(040) <= "00000000";
    -- MEMORY(041) <= "00000000";
    -- MEMORY(042) <= "00000000";
    -- MEMORY(043) <= "00000000";
    -- 
    -- MEMORY(044) <= "00000000";
    -- MEMORY(045) <= "00000000";
    -- MEMORY(046) <= "00000000";
    -- MEMORY(047) <= "00000000";
    -- 
    -- MEMORY(048) <= "00001000";
    -- MEMORY(049) <= "01100011";
    -- MEMORY(050) <= "00000000";
    -- MEMORY(051) <= "00000001";
    -- 
    -- MEMORY(052) <= "00000000";
    -- MEMORY(053) <= "00000000";
    -- MEMORY(054) <= "00000000";
    -- MEMORY(055) <= "00000000";
    -- 
    -- MEMORY(056) <= "00000000";
    -- MEMORY(057) <= "00000000";
    -- MEMORY(058) <= "00000000";
    -- MEMORY(059) <= "00000000";
    -- 
    -- MEMORY(060) <= "00000000";
    -- MEMORY(061) <= "00000000";
    -- MEMORY(062) <= "00000000";
    -- MEMORY(063) <= "00000000";
    -- 
    -- MEMORY(064) <= "00100000";
    -- MEMORY(065) <= "01100010";
    -- MEMORY(066) <= "00000000";
    -- MEMORY(067) <= "00000110";
    -- 
    -- MEMORY(068) <= "00000000";
    -- MEMORY(069) <= "00000000";
    -- MEMORY(070) <= "00000000";
    -- MEMORY(071) <= "00000000";
    -- 
    -- MEMORY(072) <= "00000000";
    -- MEMORY(073) <= "00000000";
    -- MEMORY(074) <= "00000000";
    -- MEMORY(075) <= "00000000";
    -- 
    -- MEMORY(076) <= "00000000";
    -- MEMORY(077) <= "00000000";
    -- MEMORY(078) <= "00000000";
    -- MEMORY(079) <= "00000000";
    -- 
    -- MEMORY(080) <= "00000000";
    -- MEMORY(081) <= "00000000";
    -- MEMORY(082) <= "00000000";
    -- MEMORY(083) <= "00000000";
    -- 
    -- MEMORY(084) <= "00100100";
    -- MEMORY(085) <= "00000000";
    -- MEMORY(086) <= "00000000";
    -- MEMORY(087) <= "00000111";
    -- 
    -- MEMORY(088) <= "00000000";
    -- MEMORY(089) <= "00000000";
    -- MEMORY(090) <= "00000000";
    -- MEMORY(091) <= "00000000";
    -- 
    -- MEMORY(092) <= "00000000";
    -- MEMORY(093) <= "00000000";
    -- MEMORY(094) <= "00000000";
    -- MEMORY(095) <= "00000000";
    -- 
    -- MEMORY(096) <= "00000100";
    -- MEMORY(097) <= "00100010";
    -- MEMORY(098) <= "00001000";
    -- MEMORY(099) <= "00100010";

    PROCESS (ADDRESS)
    BEGIN
        INSTRUCTION <= MEMORY(TO_INTEGER(UNSIGNED(ADDRESS))) &
            MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 1) &
            MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 2) &
            MEMORY(TO_INTEGER(UNSIGNED(ADDRESS)) + 3);
    END PROCESS;
END;